0A
1B
2C
3D
4E
5F
AA
BB
CC
DD
EE
FF
